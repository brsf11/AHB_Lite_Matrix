module ahb_lite_matrix();

endmodule