// *****************************************************************************
// (c) Copyright 2022-2032 , Inc. All rights reserved.
// Module Name  :
// Design Name  :
// Project Name :
// Create Date  : 2022-12-21
// Description  :
//
// *****************************************************************************

// -------------------------------------------------------------------
// Constant Parameter
// -------------------------------------------------------------------

// -------------------------------------------------------------------
// Internal Signals Declarations
// -------------------------------------------------------------------

// -------------------------------------------------------------------
// initial
// -------------------------------------------------------------------
`include "common/task.sv"


initial begin
  bit [31:0] rdata;
  #300;
  
  m0_test(32'h0000_0000);
  m0_test(32'h1000_0000);
  m0_test(32'h5000_0000);
end

initial begin
  bit [31:0] rdata;
  #300;
  
  m1_test(32'h0000_0010);
  m1_test(32'h2000_0000);
  m1_test(32'h6000_0000);
end

initial begin
  bit [31:0] rdata;
  #300;
  
  m2_test(32'h0000_0020);
  m2_test(32'h3000_0000);
  m2_test(32'h3000_0020);
end

initial begin
  bit [31:0] rdata;
  #300;
  
  m3_test(32'h0000_0030);
  m3_test(32'h4000_0000);
end

initial begin
  #10000;
  $finish();
end


// -------------------------------------------------------------------
// Main Code
// -------------------------------------------------------------------


// -------------------------------------------------------------------
// Assertion Declarations
// -------------------------------------------------------------------
`ifdef SOC_ASSERT_ON

`endif
